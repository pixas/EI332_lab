module sc_datamem (addr, datain, we, clock, mem_clk, dmem_clk, dataout);
 
   input  [31:0]  addr;
   input  [31:0]  datain;
   
   input          we, clock,mem_clk;
   output [31:0]  dataout;
   output         dmem_clk;
   
   wire           dmem_clk;    
   wire           write_enable; 
   assign         write_enable = we & ~clock; 
   
   assign         dmem_clk = mem_clk & ( ~ clock) ; // 分频
   
   lpm_ram_dq_dram  dram(addr[6:2], dmem_clk, datain, write_enable, dataout );

endmodule 